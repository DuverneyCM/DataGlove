library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_misc.all;
use work.spi_param.all;

entity spi_controller_fsm is
	port
	(
		-- Input ports
		ISPI_CLK			: in  std_logic;
		IRSTN				: in  std_logic;
		start				: in	std_logic;
		
		oSPI_END			: out std_logic;
		
		-- Output ports
		R_nW				: out  std_logic;
		MB					: out  std_logic;
		iAddress			: out  std_logic_vector(5 downto 0);
		iData				: out  std_logic_vector(7 downto 0);
		iSPI_GO			: out  std_logic;	
		
		oSPI_CSN			: out std_logic
	);
end spi_controller_fsm;


architecture rtl of spi_controller_fsm is

	-- Build an enumerated type for the state machine
	type state_type is (s0, s1, s2, s3);
	-- Register to hold the current state
	signal state   : state_type;

begin

	-- Logic to advance to the next state
	process (clk, reset)
	begin
		if reset = '1' then
			state <= s0;
		elsif (rising_edge(clk)) then
			case state is
				when s0=>
					if input = '1' then
						state <= s1;
					else
						state <= s0;
					end if;
				when s1=>
					if input = '1' then
						state <= s2;
					else
						state <= s1;
					end if;
				when s2=>
					if input = '1' then
						state <= s3;
					else
						state <= s2;
					end if;
				when s3 =>
					if input = '1' then
						state <= s0;
					else
						state <= s3;
					end if;
			end case;
		end if;
	end process;

	-- Output depends solely on the current state
	process (state)
	begin
		case state is
			when s0 =>
				output <= "00";
			when s1 =>
				output <= "01";
			when s2 =>
				output <= "10";
			when s3 =>
				output <= "11";
		end case;
	end process;

end rtl;
